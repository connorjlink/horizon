-- Horizon: entity.vhd
-- (c) 2026 Connor J. Link. All rights reserved.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.types.all;

entity <ENTITY_NAME> is
    port(
        i_Clock : in  std_logic;
        i_Reset : in  std_logic
    );
end <ENTITY_NAME>;

architecture implementation of <ENTITY_NAME> is
begin

    -- TODO: implementation here

end implementation;